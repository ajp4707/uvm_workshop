package cat_dog_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"  
  `include "cat.svh" 
  `include "dog.svh" 
endpackage
