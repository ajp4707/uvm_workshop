class monitor;

   // Please declare a virtual interface of type counter_if called i.

   // Please create a constructor called new that accepts a 
   // virtual interface counter_if as an argument

   // Please create a task called run that loops forever and 
   // prints the counter's out on the negative  edge of i.clk.

endclass // monitor


