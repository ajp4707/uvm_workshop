package memory_pkg;
   import uvm_pkg::*;

   virtual interface memory_if global_mif;

`include "uvm_macros.svh"
`include "quiet_test.svh"   
`include "verbose_test.svh"
endpackage: memory_pkg


