import uvm_pkg::*;
import cat_dog_pkg::*;

module top;
  
  initial run_test();
  
endmodule

