package memory_pkg;
   import uvm_pkg::*;
`include "tester.svh"
`include "monitor.svh"
`include "scoreboard.svh"
endpackage // memory_pkg
   
   
   