import uvm_pkg::*;
import producer_consumer_pkg::*;

module top;

  initial run_test("producer_consumer_test");  

endmodule: top
