package mypackage;
   integer a;
endpackage // mypackage
