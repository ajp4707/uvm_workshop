package multi_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "animal_pen.svh"
  `include "multi.svh" 
   
endpackage
