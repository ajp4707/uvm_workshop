package counter_pkg;
   // Please include tester.svh
`include "tester.svh"
   // Please include checker.svh
`include "ctr_checker.svh"
   // Please include monitor.svh
`include "monitor.svh"
endpackage // counter_pkg
   