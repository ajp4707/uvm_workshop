
module top;
   initial       $timeformat(-12, 0, " ps");
   mod1 m1();
   mod2 m2();
endmodule // top
