package counter_pkg;
   // Please include tester.svh
   // Please include ctr_checker.svh
   // Please include monitor.svh
  
endpackage // counter_pkg

